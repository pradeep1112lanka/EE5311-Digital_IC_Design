** sch_path: /home/ee22b074/ee5311/tutorial_6/test/fulladder.sch
.subckt fulladder DVDD A B Cin Cout Sum DGND
*.PININFO Cout:O Sum:O A:I B:I Cin:I DVDD:B DGND:B
XM25 net3 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM26 net3 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM27 net2 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM28 net2 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM29 net2 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM30 net2 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM31 Cout B net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM32 Cout B net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM33 Cout Cin net2 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM34 Cout Cin net2 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM35 net6 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM36 net6 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM37 net6 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM38 net6 B DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM39 net6 Cin DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM40 net6 Cin DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM41 Sum Cout net6 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM42 Sum Cout net6 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM43 net7 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM44 net7 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM45 net7 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM46 net8 B net7 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM47 net8 B net7 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM48 net8 B net7 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM49 Sum Cin net8 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM50 Sum Cin net8 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM51 Sum Cin net8 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM52 Cout A net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM53 Cout A net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM54 net1 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM55 net1 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM56 Cout Cin net4 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM57 Cout Cin net4 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM58 net4 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM59 net4 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM60 net4 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM61 net4 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM62 Sum Cout net5 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM63 Sum Cout net5 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM64 net5 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM65 net5 A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM66 net5 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM67 net5 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM68 net5 Cin DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM69 net5 Cin DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM70 Sum Cin net9 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM71 Sum Cin net9 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM72 net9 A net10 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM73 net9 A net10 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM74 net10 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM75 net10 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM76 Sum Cin net9 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM77 net9 A net10 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM78 net10 B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.GLOBAL GND
.end
