* NGSPICE file created from TOP.ext - technology: sky130A

.subckt TOP B1 S1 A1 A0 B0 S0 B2 S2 A2 B3 S3 A3 B4 S4 A4 B5 S5 A5 B6 S6 A6 B7 S7 A7
+ DVDD DGND C7
X0 a_1406_n143# B0 a_1136_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X1 DVDD A7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_414_n6526# B7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X3 S1 C7 a_1403_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X4 a_1403_n1032# B1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X5 a_n670_n412# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X6 a_n313_n2133# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X7 a_416_n412# C7 S0 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X8 DGND B0 a_n310_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X9 a_413_n1301# B1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X10 DVDD A1 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X11 a_n672_n6257# A7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X12 S0 C7 a_1406_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X13 S6 C7 a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X14 a_1134_n2716# A3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X15 S3 C7 a_1404_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X16 a_413_n5405# C7 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X17 a_414_n2716# A3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X18 DGND A4 a_n312_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X19 a_414_n2985# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X20 a_1133_n2133# B2 a_1403_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X21 a_416_n143# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X22 DVDD A3 a_n672_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X23 DGND A6 a_1133_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X24 DVDD B6 a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X25 a_413_n2133# C7 S2 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X26 DGND B3 a_n312_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X27 a_n312_n3687# C7 C7 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X28 C7 C7 a_n312_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X29 S0 C7 a_1406_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X30 a_1134_n2716# A3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X31 DGND A0 a_416_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X32 a_n313_n5405# C7 C7 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X33 a_n673_n5674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X34 DGND A7 a_n312_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X35 DGND C7 a_413_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X36 a_1404_n3956# C7 S4 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X37 S4 C7 a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X38 S0 C7 a_416_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X39 a_n312_n6257# C7 a_n582_n6526# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X40 a_n582_n6526# C7 a_n312_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X41 DGND B4 a_414_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X42 a_414_n3687# B4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X43 a_1133_n5405# A6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X44 a_1406_n143# C7 S0 DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X45 S6 C7 a_1403_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X46 a_1134_n2985# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X47 a_413_n5405# A6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X48 a_413_n5674# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X49 a_416_n412# B0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X50 a_414_n2985# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X51 a_n673_n1032# B1 C7 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X52 C7 B1 a_n673_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X53 S5 C7 a_1405_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X54 a_1405_n4539# B5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X55 DGND A3 a_n672_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X56 DGND B6 a_n313_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X57 a_415_n4808# B5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X58 DVDD A5 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X59 a_1133_n1864# B2 a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X60 a_1133_n5405# A6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X61 S7 C7 a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X62 DGND A5 a_n671_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X63 a_1404_n6526# C7 S7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X64 a_1134_n2985# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X65 a_413_n1864# C7 S2 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X66 a_414_n6257# B7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X67 DGND B7 a_414_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X68 a_n670_n143# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X69 a_1403_n1301# C7 S1 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X70 S1 C7 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X71 a_416_n143# C7 S0 DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X72 DGND A2 a_n673_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X73 DVDD B0 a_n310_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X74 a_413_n1032# B1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X75 DGND B1 a_413_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X76 a_n313_n5674# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X77 S0 C7 a_1406_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X78 a_1404_n2716# B3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X79 a_n312_n2716# B3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X80 DGND B0 a_416_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X81 DGND A0 a_n310_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X82 DVDD A4 a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X83 S3 C7 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X84 DGND A4 a_1134_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X85 a_1403_n2133# B2 a_1133_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X86 a_n672_n2716# B3 C7 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X87 a_1133_n5674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X88 DGND A2 a_413_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X89 DVDD A6 a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X90 C7 C7 a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X91 a_413_n5674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X92 a_n312_n3956# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X93 DVDD A0 a_416_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X94 DGND C7 a_414_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X95 C7 C7 a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X96 DVDD A7 a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X97 a_416_n412# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X98 a_1133_n5674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X99 DGND A7 a_1134_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X100 DGND A1 a_1133_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X101 S4 C7 a_1404_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X102 a_1404_n3687# C7 S4 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X103 a_n582_n6526# C7 a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X104 a_n312_n6526# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X105 DVDD B4 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X106 a_414_n3956# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X107 a_n313_n5405# B6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X108 DVDD A2 a_n673_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X109 a_1403_n5405# B6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X110 DGND C7 a_416_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X111 a_1404_n2985# B3 a_1134_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X112 a_n312_n2985# B3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X113 a_416_n143# B0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X114 S6 C7 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X115 DGND C7 a_414_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X116 S3 C7 a_414_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X117 C7 B1 a_n673_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X118 DGND B4 a_n312_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X119 a_n673_n1301# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X120 DGND C7 a_413_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X121 S5 C7 a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X122 a_1405_n4808# C7 S5 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X123 a_n672_n2985# B3 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X124 a_415_n4539# B5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X125 DGND B5 a_415_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X126 a_1403_n1864# B2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X127 DGND A6 a_n313_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X128 DVDD A5 a_n671_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X129 a_1404_n6257# C7 S7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X130 a_n671_n4808# B5 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X131 S7 C7 a_1404_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X132 DVDD A2 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X133 DVDD B7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X134 a_414_n6526# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X135 a_1403_n1032# C7 S1 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X136 S1 C7 a_1403_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X137 a_n673_n2133# B2 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X138 DVDD B1 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X139 C7 C7 a_n313_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X140 a_413_n1301# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X141 a_1136_n412# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X142 DGND B7 a_n312_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X143 DVDD B0 a_416_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X144 a_1134_n2716# B3 a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X145 DVDD A0 a_n310_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X146 DGND B1 a_n313_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X147 a_414_n2716# C7 S3 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X148 a_1134_n3956# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X149 DVDD A4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X150 a_414_n3956# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X151 S2 C7 a_1403_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X152 a_n313_n5674# B6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X153 C7 B3 a_n672_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X154 a_1403_n5674# B6 a_1133_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X155 a_413_n2133# B2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X156 S6 C7 a_413_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X157 DGND A4 a_n672_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X158 a_n313_n1301# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X159 DVDD C7 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X160 DGND A5 a_1135_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X161 a_1134_n3956# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X162 a_416_n143# C7 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X163 DVDD A7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X164 a_1134_n6526# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X165 a_414_n6526# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X166 DVDD A1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X167 a_1133_n1301# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X168 S4 C7 a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X169 a_413_n1301# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X170 DGND A7 a_n672_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X171 DGND C7 a_415_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X172 a_414_n3687# C7 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X173 DVDD C7 a_416_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X174 a_n673_n1864# B2 C7 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X175 a_1133_n5405# B6 a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X176 a_n310_n412# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X177 a_1134_n2985# B3 a_1404_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X178 DVDD C7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X179 a_413_n5405# C7 S6 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X180 a_1134_n6526# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X181 DVDD B4 a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X182 a_414_n2985# C7 S3 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X183 a_n673_n1032# A1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X184 DVDD C7 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X185 a_1133_n1301# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X186 a_1405_n4539# C7 S5 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X187 S5 C7 a_1405_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X188 C7 B3 a_n672_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X189 DVDD B5 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X190 a_415_n4808# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X191 S2 C7 a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X192 C7 B5 a_n671_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X193 a_n671_n4539# B5 C7 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X194 S7 C7 a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X195 a_413_n1864# B2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X196 a_414_n6257# C7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X197 S1 C7 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X198 DGND B5 a_n311_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X199 C7 B2 a_n673_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X200 a_1136_n143# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X201 a_413_n1032# C7 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X202 a_n313_n5674# A6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X203 C7 C7 a_n310_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X204 DVDD B7 a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X205 a_1404_n2716# B3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X206 DVDD B1 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X207 a_n312_n3956# B4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X208 a_1134_n3687# A4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X209 DVDD A3 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X210 a_1404_n3956# B4 a_1134_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X211 DGND A1 a_n313_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X212 a_414_n3687# A4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X213 a_1403_n2133# C7 S2 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X214 S4 C7 a_414_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X215 a_n672_n2716# A3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X216 a_1133_n5674# B6 a_1403_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X217 DGND B2 a_413_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X218 a_n672_n3956# B4 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X219 DVDD A4 a_n672_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X220 a_413_n5674# C7 S6 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X221 C7 C7 a_n313_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X222 a_n313_n1032# C7 C7 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X223 DVDD A5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X224 a_1134_n3687# A4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X225 a_1135_n4808# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X226 a_n310_n412# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X227 DVDD A6 a_n673_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X228 a_415_n4808# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X229 a_1134_n6257# A7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X230 a_n312_n6526# B7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X231 a_1404_n6526# B7 a_1134_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X232 a_414_n6257# A7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X233 S7 a_n582_n6526# a_414_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X234 a_n313_n1301# B1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X235 a_1133_n1032# A1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X236 a_1403_n1301# B1 a_1133_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X237 a_413_n1032# A1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X238 DVDD A7 a_n672_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X239 S1 C7 a_413_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X240 a_n672_n6526# B7 a_n582_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X241 DVDD C7 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X242 a_1135_n4808# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X243 C7 B2 a_n673_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X244 a_1403_n5405# B6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X245 a_1404_n2985# B3 a_1134_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X246 a_1134_n6257# A7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X247 DVDD A6 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X248 DGND A3 a_414_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X249 a_1133_n1032# A1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X250 DGND A2 a_1133_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X251 DGND A0 a_n670_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X252 S5 C7 a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X253 a_n312_n2716# C7 C7 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X254 a_n672_n2985# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X255 a_415_n4539# C7 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X256 a_1403_n1864# C7 S2 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X257 a_n671_n4808# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X258 C7 B5 a_n671_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X259 DVDD B2 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X260 DVDD B5 a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X261 a_n673_n2133# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X262 a_n310_n412# B0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X263 DGND C7 a_413_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X264 DGND A6 a_n673_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X265 C7 C7 a_n310_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.123 pd=1.12 as=0.084 ps=0.76 w=1.66 l=0.15
X266 DGND A0 a_1136_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X267 S3 C7 a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X268 a_1404_n3687# B4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X269 a_n312_n3687# B4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X270 a_414_n2716# B3 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X271 a_n670_n412# B0 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X272 a_1134_n3956# B4 a_1404_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X273 DVDD A1 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X274 S4 C7 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X275 S2 C7 a_1403_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X276 a_414_n3956# C7 S4 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X277 a_1403_n5674# B6 a_1133_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X278 a_413_n2133# C7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X279 DGND A6 a_413_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X280 C7 B4 a_n672_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X281 a_n672_n3687# B4 C7 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X282 a_n313_n1301# A1 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X283 C7 C7 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X284 DGND B2 a_n313_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X285 a_n311_n4808# B5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X286 a_1135_n4539# A5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X287 a_1405_n4808# B5 a_1135_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X288 a_n312_n2985# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X289 a_1136_n412# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X290 a_n673_n5405# B6 C7 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X291 a_415_n4539# A5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X292 S5 C7 a_415_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X293 DVDD A2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X294 a_n312_n6257# B7 DVDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X295 a_n311_n4808# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X296 a_1404_n6257# B7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X297 a_1134_n6526# B7 a_1404_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X298 S7 a_n582_n6526# a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X299 a_414_n6526# a_n582_n6526# S7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X300 a_n313_n1032# B1 DVDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X301 C7 B0 a_n670_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X302 a_1403_n1032# B1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X303 a_1133_n1301# B1 a_1403_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X304 a_n313_n2133# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X305 S1 C7 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X306 a_n672_n6257# B7 a_n582_n6526# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X307 a_413_n1301# C7 S1 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X308 a_n582_n6526# B7 a_n672_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X309 a_1135_n4539# A5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X310 a_n673_n1864# A2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X311 S6 C7 a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X312 DVDD A3 a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X313 DVDD C7 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X314 S3 C7 a_1404_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X315 a_413_n5405# B6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X316 a_414_n2985# B3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X317 DVDD A0 a_n670_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X318 a_1133_n2133# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X319 a_1406_n412# B0 a_1136_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X320 C7 C7 a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X321 a_413_n2133# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X322 a_n671_n4539# A5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X323 S2 C7 a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X324 a_413_n1864# C7 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X325 a_n310_n143# B0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X326 a_1133_n2133# A2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X327 a_n673_n5674# B6 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X328 DVDD B2 a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X329 DVDD A0 a_1136_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X330 a_1404_n2716# C7 S3 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X331 a_n670_n143# B0 C7 DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X332 a_1134_n3687# B4 a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X333 DVDD B3 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X334 a_1136_n412# B0 a_1406_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X335 a_1404_n3956# B4 a_1134_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X336 a_414_n3687# C7 S4 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X337 DGND A4 a_414_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X338 a_n313_n1864# C7 C7 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X339 S6 C7 a_1403_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X340 DGND A3 a_n312_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X341 C7 B4 a_n672_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X342 a_413_n5674# B6 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X343 a_n672_n3956# A4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X344 DGND A5 a_n311_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X345 DGND A1 a_n673_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X346 a_n311_n4539# B5 DVDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X347 a_1405_n4539# B5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X348 a_1136_n143# A0 DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X349 a_1135_n4808# B5 a_1405_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X350 C7 C7 a_n312_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X351 DGND A2 a_n313_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X352 C7 B6 a_n673_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X353 S5 C7 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X354 a_415_n4808# C7 S5 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X355 a_n311_n4539# C7 C7 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X356 a_1133_n1864# A2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X357 C7 C7 a_n311_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X358 a_1134_n6257# B7 a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X359 a_1404_n6526# B7 a_1134_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X360 a_413_n1864# A2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X361 C7 B0 a_n670_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X362 a_414_n6257# a_n582_n6526# S7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X363 DGND A7 a_414_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X364 a_1406_n412# B0 a_1136_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X365 a_1133_n1032# B1 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X366 a_1403_n1301# B1 a_1133_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X367 C7 C7 a_n313_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X368 DGND A1 a_413_n1301# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X369 a_413_n1032# C7 S1 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X370 a_n582_n6526# B7 a_n672_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X371 a_n672_n6526# A7 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X372 a_1403_n5405# C7 S6 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X373 DVDD A3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X374 a_1133_n1864# A2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X375 a_1404_n2985# C7 S3 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X376 DVDD B6 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X377 DGND B3 a_414_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X378 a_1406_n143# B0 a_1136_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X379 a_n313_n2133# B2 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X380 a_1403_n2133# B2 a_1133_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X381 a_416_n412# A0 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X382 S2 C7 a_413_n2133# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X383 a_n312_n3956# C7 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X384 S0 C7 a_1406_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X385 DVDD C7 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X386 C7 B6 a_n673_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X387 DVDD A2 a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X388 S3 C7 a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X389 a_1136_n143# B0 a_1406_n143# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X390 a_414_n2716# C7 DVDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X391 a_1404_n3687# B4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X392 S4 C7 a_1404_n3956# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X393 S0 C7 a_416_n412# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X394 a_n312_n6526# C7 a_n582_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X395 DVDD A4 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X396 a_414_n3956# B4 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X397 C7 C7 a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X398 DVDD A6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X399 a_1403_n5674# C7 S6 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X400 DGND A3 a_1134_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X401 DVDD B3 a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X402 a_1406_n412# C7 S0 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X403 a_n672_n3687# A4 DVDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X404 DGND B6 a_413_n5674# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X405 DVDD A5 a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X406 DVDD A1 a_n673_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X407 a_n673_n1301# B1 C7 DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X408 a_1135_n4539# B5 a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X409 a_1405_n4808# B5 a_1135_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X410 a_n312_n2985# A3 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X411 a_n673_n5405# A6 DVDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X412 DGND A5 a_415_n4808# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X413 a_415_n4539# C7 S5 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X414 a_n313_n1864# B2 DVDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X415 C7 C7 a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X416 a_1403_n1864# B2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X417 DVDD C7 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X418 a_1404_n6257# B7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X419 a_n311_n4808# A5 DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X420 S7 C7 a_1404_n6526# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X421 DGND C7 a_414_n2985# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X422 S2 C7 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
.ends

