* NGSPICE file created from rippleadder.ext - technology: sky130A

.subckt rippleadder A7 B7 A6 B6 A5 A4 A3 A2 A1 S1 S2 S3 S4 S5 S6 S7 A0 DGNDD DVDDD
+ B1 B0 C0 S0 B2 B3 B4 B5 C7
X0 a_1406_n143# B0 a_1136_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X1 DVDDD A7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X2 a_414_n6526# B7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X3 S1 C0 a_1403_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X4 a_1403_n1032# B1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X5 a_n670_n412# A0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X6 a_n313_n2133# A2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X7 a_416_n412# C0 S0 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X8 DGNDD B0 a_n310_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X9 a_413_n1301# B1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X10 DVDDD A1 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X11 a_n672_n6257# A7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X12 S0 a_n250_n452# a_1406_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X13 S6 a_n581_n4808# a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X14 a_1134_n2716# A3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X15 S3 a_n583_n2133# a_1404_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X16 a_413_n5405# a_n581_n4808# DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X17 a_414_n2716# A3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X18 DGNDD A4 a_n312_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X19 a_414_n2985# a_n583_n2133# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X20 a_1133_n2133# B2 a_1403_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X21 a_416_n143# A0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X22 DVDDD A3 a_n672_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X23 DGNDD A6 a_1133_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X24 DVDDD B6 a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X25 a_413_n2133# a_n583_n2133# S2 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X26 DGNDD B3 a_n312_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X27 a_n312_n3687# a_n582_n2985# a_n582_n3956# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X28 a_n582_n3956# a_n582_n2985# a_n312_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X29 S0 a_n250_n452# a_1406_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X30 a_1134_n2716# A3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X31 DGNDD A0 a_416_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X32 a_n313_n5405# a_n581_n4808# a_n583_n5674# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X33 a_n673_n5674# A6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X34 DGNDD A7 a_n312_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X35 DGNDD a_n581_n4808# a_413_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X36 a_1404_n3956# a_n582_n2985# S4 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X37 S4 a_n582_n2985# a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X38 S0 C0 a_416_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X39 a_n312_n6257# a_n583_n5674# C7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X40 C7 a_n583_n5674# a_n312_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X41 DGNDD B4 a_414_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X42 a_414_n3687# B4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X43 a_1133_n5405# A6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X44 a_1406_n143# a_n250_n452# S0 DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X45 S6 a_n581_n4808# a_1403_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X46 a_1134_n2985# A3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X47 a_413_n5405# A6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X48 a_413_n5674# a_n581_n4808# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X49 a_416_n412# B0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X50 a_414_n2985# A3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X51 a_n673_n1032# B1 a_n583_n1301# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X52 a_n583_n1301# B1 a_n673_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X53 S5 a_n582_n3956# a_1405_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X54 a_1405_n4539# B5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X55 DGNDD A3 a_n672_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X56 DGNDD B6 a_n313_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X57 a_415_n4808# B5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X58 DVDDD A5 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X59 a_1133_n1864# B2 a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X60 a_1133_n5405# A6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X61 S7 a_n583_n5674# a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X62 DGNDD A5 a_n671_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X63 a_1404_n6526# a_n583_n5674# S7 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X64 a_1134_n2985# A3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X65 a_413_n1864# a_n583_n2133# S2 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X66 a_414_n6257# B7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X67 DGNDD B7 a_414_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X68 a_n670_n143# A0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X69 a_1403_n1301# C0 S1 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X70 S1 C0 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X71 a_416_n143# C0 S0 DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X72 DGNDD A2 a_n673_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X73 DVDDD B0 a_n310_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X74 a_413_n1032# B1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X75 DGNDD B1 a_413_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X76 a_n313_n5674# a_n581_n4808# a_n583_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X77 S0 a_n250_n452# a_1406_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X78 a_1404_n2716# B3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X79 a_n312_n2716# B3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X80 DGNDD B0 a_416_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X81 DGNDD A0 a_n310_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X82 DVDDD A4 a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X83 S3 a_n582_n2985# a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X84 DGNDD A4 a_1134_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X85 a_1403_n2133# B2 a_1133_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X86 a_n672_n2716# B3 a_n582_n2985# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X87 a_1133_n5674# A6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X88 DGNDD A2 a_413_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X89 DVDDD A6 a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X90 a_n582_n3956# a_n582_n2985# a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X91 a_413_n5674# A6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X92 a_n312_n3956# A4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X93 DVDDD A0 a_416_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X94 DGNDD a_n582_n2985# a_414_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X95 a_n583_n5674# a_n581_n4808# a_n313_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X96 DVDDD A7 a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X97 a_416_n412# a_n250_n452# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X98 a_1133_n5674# A6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X99 DGNDD A7 a_1134_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X100 DGNDD A1 a_1133_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X101 S4 a_n582_n2985# a_1404_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X102 a_1404_n3687# a_n582_n2985# S4 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X103 C7 a_n583_n5674# a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X104 a_n312_n6526# A7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X105 DVDDD B4 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X106 a_414_n3956# a_n582_n2985# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X107 a_n313_n5405# B6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X108 DVDDD A2 a_n673_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X109 a_1403_n5405# B6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X110 DGNDD a_n250_n452# a_416_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X111 a_1404_n2985# B3 a_1134_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X112 a_n312_n2985# B3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X113 a_416_n143# B0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X114 S6 a_n583_n5674# a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X115 DGNDD a_n583_n5674# a_414_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X116 S3 a_n582_n2985# a_414_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X117 a_n583_n1301# B1 a_n673_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X118 DGNDD B4 a_n312_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X119 a_n673_n1301# A1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X120 DGNDD C0 a_413_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X121 S5 a_n582_n3956# a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X122 a_1405_n4808# a_n582_n3956# S5 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X123 a_n672_n2985# B3 a_n582_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X124 a_415_n4539# B5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X125 DGNDD B5 a_415_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X126 a_1403_n1864# B2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X127 DGNDD A6 a_n313_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X128 DVDDD A5 a_n671_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X129 a_1404_n6257# a_n583_n5674# S7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X130 a_n671_n4808# B5 a_n581_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X131 S7 a_n583_n5674# a_1404_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X132 DVDDD A2 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X133 DVDDD B7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X134 a_414_n6526# a_n583_n5674# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X135 a_1403_n1032# C0 S1 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X136 S1 C0 a_1403_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X137 a_n673_n2133# B2 a_n583_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X138 DVDDD B1 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X139 a_n583_n5674# a_n581_n4808# a_n313_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X140 a_413_n1301# C0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X141 a_1136_n412# A0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X142 DGNDD B7 a_n312_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X143 DVDDD B0 a_416_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X144 a_1134_n2716# B3 a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X145 DVDDD A0 a_n310_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X146 DGNDD B1 a_n313_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X147 a_414_n2716# a_n582_n2985# S3 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X148 a_1134_n3956# A4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X149 DVDDD A4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X150 a_414_n3956# A4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X151 S2 a_n583_n1301# a_1403_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X152 a_n313_n5674# B6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X153 a_n582_n2985# B3 a_n672_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X154 a_1403_n5674# B6 a_1133_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X155 a_413_n2133# B2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X156 S6 a_n583_n5674# a_413_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X157 DGNDD A4 a_n672_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X158 a_n313_n1301# C0 a_n583_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X159 DVDDD a_n582_n2985# a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X160 DGNDD A5 a_1135_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X161 a_1134_n3956# A4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X162 a_416_n143# a_n250_n452# DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X163 DVDDD A7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X164 a_1134_n6526# A7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X165 a_414_n6526# A7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X166 DVDDD A1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X167 a_1133_n1301# A1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X168 S4 a_n582_n2985# a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X169 a_413_n1301# A1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X170 DGNDD A7 a_n672_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X171 DGNDD a_n582_n3956# a_415_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X172 a_414_n3687# a_n582_n2985# DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X173 DVDDD a_n250_n452# a_416_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X174 a_n673_n1864# B2 a_n583_n2133# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X175 a_1133_n5405# B6 a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X176 a_n310_n412# a_n250_n452# C0 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X177 a_1134_n2985# B3 a_1404_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X178 DVDDD a_n583_n5674# a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X179 a_413_n5405# a_n583_n5674# S6 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X180 a_1134_n6526# A7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X181 DVDDD B4 a_n312_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X182 a_414_n2985# a_n582_n2985# S3 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X183 a_n673_n1032# A1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X184 DVDDD C0 a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X185 a_1133_n1301# A1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X186 a_1405_n4539# a_n582_n3956# S5 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X187 S5 a_n582_n3956# a_1405_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X188 a_n582_n2985# B3 a_n672_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X189 DVDDD B5 a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X190 a_415_n4808# a_n582_n3956# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X191 S2 a_n583_n1301# a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X192 a_n581_n4808# B5 a_n671_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X193 a_n671_n4539# B5 a_n581_n4808# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X194 S7 a_n583_n5674# a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X195 a_413_n1864# B2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X196 a_414_n6257# a_n583_n5674# DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X197 S1 C0 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X198 DGNDD B5 a_n311_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X199 a_n583_n2133# B2 a_n673_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X200 a_1136_n143# A0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X201 a_413_n1032# C0 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X202 a_n313_n5674# A6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X203 C0 a_n250_n452# a_n310_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X204 DVDDD B7 a_n312_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X205 a_1404_n2716# B3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X206 DVDDD B1 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X207 a_n312_n3956# B4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X208 a_1134_n3687# A4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X209 DVDDD A3 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X210 a_1404_n3956# B4 a_1134_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X211 DGNDD A1 a_n313_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X212 a_414_n3687# A4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X213 a_1403_n2133# a_n583_n1301# S2 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X214 S4 a_n582_n3956# a_414_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X215 a_n672_n2716# A3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X216 a_1133_n5674# B6 a_1403_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X217 DGNDD B2 a_413_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X218 a_n672_n3956# B4 a_n582_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X219 DVDDD A4 a_n672_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X220 a_413_n5674# a_n583_n5674# S6 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X221 a_n583_n1301# C0 a_n313_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X222 a_n313_n1032# C0 a_n583_n1301# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X223 DVDDD A5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X224 a_1134_n3687# A4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X225 a_1135_n4808# A5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X226 a_n310_n412# A0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X227 DVDDD A6 a_n673_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X228 a_415_n4808# A5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X229 a_1134_n6257# A7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X230 a_n312_n6526# B7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X231 a_1404_n6526# B7 a_1134_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X232 a_414_n6257# A7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X233 S7 C7 a_414_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X234 a_n313_n1301# B1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X235 a_1133_n1032# A1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X236 a_1403_n1301# B1 a_1133_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X237 a_413_n1032# A1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X238 DVDDD A7 a_n672_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X239 S1 a_n583_n1301# a_413_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X240 a_n672_n6526# B7 C7 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X241 DVDDD a_n582_n3956# a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X242 a_1135_n4808# A5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X243 a_n583_n2133# B2 a_n673_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X244 a_1403_n5405# B6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X245 a_1404_n2985# B3 a_1134_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X246 a_1134_n6257# A7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X247 DVDDD A6 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X248 DGNDD A3 a_414_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X249 a_1133_n1032# A1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X250 DGNDD A2 a_1133_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X251 DGNDD A0 a_n670_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X252 S5 a_n582_n3956# a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X253 a_n312_n2716# a_n583_n2133# a_n582_n2985# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X254 a_n672_n2985# A3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X255 a_415_n4539# a_n582_n3956# DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X256 a_1403_n1864# a_n583_n1301# S2 w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X257 a_n671_n4808# A5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X258 a_n581_n4808# B5 a_n671_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X259 DVDDD B2 a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X260 DVDDD B5 a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X261 a_n673_n2133# A2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X262 a_n310_n412# B0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X263 DGNDD a_n583_n1301# a_413_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X264 DGNDD A6 a_n673_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X265 C0 a_n250_n452# a_n310_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.123 pd=1.12 as=0.084 ps=0.76 w=1.66 l=0.15
X266 DGNDD A0 a_1136_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X267 S3 a_n583_n2133# a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X268 a_1404_n3687# B4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X269 a_n312_n3687# B4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X270 a_414_n2716# B3 DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X271 a_n670_n412# B0 C0 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X272 a_1134_n3956# B4 a_1404_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X273 DVDDD A1 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X274 S4 a_n582_n3956# a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X275 S2 a_n583_n1301# a_1403_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X276 a_414_n3956# a_n582_n3956# S4 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X277 a_1403_n5674# B6 a_1133_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X278 a_413_n2133# a_n583_n1301# DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X279 DGNDD A6 a_413_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X280 a_n582_n3956# B4 a_n672_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X281 a_n672_n3687# B4 a_n582_n3956# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X282 a_n313_n1301# A1 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X283 a_n583_n1301# C0 a_n313_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X284 DGNDD B2 a_n313_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.063 ps=0.72 w=0.42 l=0.15
X285 a_n311_n4808# B5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X286 a_1135_n4539# A5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X287 a_1405_n4808# B5 a_1135_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X288 a_n312_n2985# a_n583_n2133# a_n582_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X289 a_1136_n412# A0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X290 a_n673_n5405# B6 a_n583_n5674# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X291 a_415_n4539# A5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X292 S5 a_n581_n4808# a_415_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X293 DVDDD A2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X294 a_n312_n6257# B7 DVDDD w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X295 a_n311_n4808# a_n582_n3956# a_n581_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X296 a_1404_n6257# B7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X297 a_1134_n6526# B7 a_1404_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X298 S7 C7 a_414_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X299 a_414_n6526# C7 S7 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X300 a_n313_n1032# B1 DVDDD w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X301 C0 B0 a_n670_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X302 a_1403_n1032# B1 a_1133_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X303 a_1133_n1301# B1 a_1403_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X304 a_n313_n2133# a_n583_n1301# a_n583_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X305 S1 a_n583_n1301# a_413_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X306 a_n672_n6257# B7 C7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X307 a_413_n1301# a_n583_n1301# S1 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X308 C7 B7 a_n672_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X309 a_1135_n4539# A5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X310 a_n673_n1864# A2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X311 S6 a_n581_n4808# a_1403_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X312 DVDDD A3 a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X313 DVDDD a_n583_n1301# a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X314 S3 a_n583_n2133# a_1404_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X315 a_413_n5405# B6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X316 a_414_n2985# B3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X317 DVDDD A0 a_n670_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X318 a_1133_n2133# A2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X319 a_1406_n412# B0 a_1136_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X320 a_n582_n2985# a_n583_n2133# a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X321 a_413_n2133# A2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X322 a_n671_n4539# A5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X323 S2 a_n583_n1301# a_1403_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X324 a_413_n1864# a_n583_n1301# DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X325 a_n310_n143# B0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X326 a_1133_n2133# A2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X327 a_n673_n5674# B6 a_n583_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X328 DVDDD B2 a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X329 DVDDD A0 a_1136_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X330 a_1404_n2716# a_n583_n2133# S3 w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X331 a_n670_n143# B0 C0 DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X332 a_1134_n3687# B4 a_1404_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X333 DVDDD B3 a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X334 a_1136_n412# B0 a_1406_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X335 a_1404_n3956# B4 a_1134_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X336 a_414_n3687# a_n582_n3956# S4 w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X337 DGNDD A4 a_414_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X338 a_n313_n1864# a_n583_n1301# a_n583_n2133# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X339 S6 a_n581_n4808# a_1403_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X340 DGNDD A3 a_n312_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X341 a_n582_n3956# B4 a_n672_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X342 a_413_n5674# B6 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X343 a_n672_n3956# A4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X344 DGNDD A5 a_n311_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X345 DGNDD A1 a_n673_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X346 a_n311_n4539# B5 DVDDD w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X347 a_1405_n4539# B5 a_1135_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X348 a_1136_n143# A0 DVDDD DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X349 a_1135_n4808# B5 a_1405_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X350 a_n582_n2985# a_n583_n2133# a_n312_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X351 DGNDD A2 a_n313_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X352 a_n583_n5674# B6 a_n673_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X353 S5 a_n581_n4808# a_415_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X354 a_415_n4808# a_n581_n4808# S5 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X355 a_n311_n4539# a_n582_n3956# a_n581_n4808# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X356 a_1133_n1864# A2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X357 a_n581_n4808# a_n582_n3956# a_n311_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X358 a_1134_n6257# B7 a_1404_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X359 a_1404_n6526# B7 a_1134_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X360 a_413_n1864# A2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X361 C0 B0 a_n670_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X362 a_414_n6257# C7 S7 w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X363 DGNDD A7 a_414_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X364 a_1406_n412# B0 a_1136_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X365 a_1133_n1032# B1 a_1403_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X366 a_1403_n1301# B1 a_1133_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X367 a_n583_n2133# a_n583_n1301# a_n313_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X368 DGNDD A1 a_413_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X369 a_413_n1032# a_n583_n1301# S1 w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X370 C7 B7 a_n672_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X371 a_n672_n6526# A7 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X372 a_1403_n5405# a_n581_n4808# S6 w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X373 DVDDD A3 a_1134_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X374 a_1133_n1864# A2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X375 a_1404_n2985# a_n583_n2133# S3 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X376 DVDDD B6 a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X377 DGNDD B3 a_414_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X378 a_1406_n143# B0 a_1136_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X379 a_n313_n2133# B2 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X380 a_1403_n2133# B2 a_1133_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X381 a_416_n412# A0 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X382 S2 a_n583_n2133# a_413_n2133# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X383 a_n312_n3956# a_n582_n2985# a_n582_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X384 S0 a_n250_n452# a_1406_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X385 DVDDD a_n583_n2133# a_414_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X386 a_n583_n5674# B6 a_n673_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X387 DVDDD A2 a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X388 S3 a_n583_n2133# a_1404_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X389 a_1136_n143# B0 a_1406_n143# DVDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X390 a_414_n2716# a_n583_n2133# DVDDD w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X391 a_1404_n3687# B4 a_1134_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X392 S4 a_n582_n2985# a_1404_n3956# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X393 S0 C0 a_416_n412# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X394 a_n312_n6526# a_n583_n5674# C7 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X395 DVDDD A4 a_414_n3687# w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X396 a_414_n3956# B4 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X397 a_n583_n2133# a_n583_n1301# a_n313_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X398 DVDDD A6 a_1133_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X399 a_1403_n5674# a_n581_n4808# S6 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X400 DGNDD A3 a_1134_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X401 DVDDD B3 a_n312_n2716# w_n825_n2794# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.126 ps=1.14 w=0.84 l=0.15
X402 a_1406_n412# a_n250_n452# S0 DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X403 a_n672_n3687# A4 DVDDD w_n825_n3765# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X404 DGNDD B6 a_413_n5674# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X405 DVDDD A5 a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X406 DVDDD A1 a_n673_n1032# w_n826_n1110# sky130_fd_pr__pfet_01v8 ad=0.12375 pd=1.125 as=0.084 ps=0.76 w=0.83 l=0.15
X407 a_n673_n1301# B1 a_n583_n1301# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X408 a_1135_n4539# B5 a_1405_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X409 a_1405_n4808# B5 a_1135_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X410 a_n312_n2985# A3 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X411 a_n673_n5405# A6 DVDDD w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X412 DGNDD A5 a_415_n4808# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X413 a_415_n4539# a_n581_n4808# S5 w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X414 a_n313_n1864# B2 DVDDD w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X415 a_n581_n4808# a_n582_n3956# a_n311_n4539# w_n824_n4617# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X416 a_1403_n1864# B2 a_1133_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X417 DVDDD a_n581_n4808# a_413_n5405# w_n826_n5483# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X418 a_1404_n6257# B7 a_1134_n6257# w_n825_n6335# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X419 a_n311_n4808# A5 DGNDD DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X420 S7 a_n583_n5674# a_1404_n6526# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X421 DGNDD a_n583_n2133# a_414_n2985# DGNDD sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X422 S2 a_n583_n2133# a_413_n1864# w_n826_n1942# sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
.ends

